

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
entity ascii2led is
Port ( ASCII : in STD_LOGIC_VECTOR (7 downto 0);
LED : out STD_LOGIC_VECTOR (6 downto 0));
end ascii2led;
architecture Behavioral of ascii2led is
--ASCII-to-seven-segment decoder
-- ASCII: in STD_LOGIC_VECTOR (7 downto 0);
-- LED: out STD_LOGIC_VECTOR (6 downto 0);
--
-- 0
-- ---
-- 5 | | 1
-- --- <- 6
-- 4 | | 2
-- ---
-- 3

BEGIN
WITH ASCII SELECT
LED <= "1000000" WHEN "00110000", --0
"1111001" WHEN "00110001", --1
"0100100" WHEN "00110010", --2
"0110000" WHEN "00110011", --3
"0011001" WHEN "00110100", --4
"0010010" WHEN "00110101", --5
"0000010" WHEN "00110110", --6
"1111000" WHEN "00110111", --7
"0000000" WHEN "00111000", --8
"0010000" WHEN "00111001", --9
"0001000" WHEN "01000001", --A
"0000011" WHEN "01000010", --B
"1000110" WHEN "01000011", --C
"0100001" WHEN "01000100", --D
"0000110" WHEN "01000101", --E
"0001110" WHEN "01000110", --F
"1000010" WHEN "01000111", --G
"0001011" WHEN "01001000", --H
"1111011" WHEN "01001001", --I
"1100001" WHEN "01001010", --J
"0001010" WHEN "01001011", --K
"1000111" WHEN "01001100", --L
"1001000" WHEN "01001101", --M
"0101011" WHEN "01001110", --N
"0100011" WHEN "01001111", --O
"0001100" WHEN "01010000", --P
"0011000" WHEN "01010001", --Q
"0101111" WHEN "01010010", --R
"0010011" WHEN "01010011", --S
"0000111" WHEN "01010100", --T
"1100011" WHEN "01010101", --U
"1000001" WHEN "01010110", --V
"0000001" WHEN "01010111", --W
"0001001" WHEN "01011000", --X
"0010001" WHEN "01011001", --Y
"1100100" WHEN "01011010", --Z
"0110110" WHEN OTHERS; -- UNDEFINED
end Behavioral;

